library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.alu_pkg.all;


architecture struct of parser_top is 

begin
     
     ---parser_logic_instance
     
     alu_top_inst : alu_top
	generic
	(
	    RESET_VALUE =>
	);
	port
	(
		sys_clk	=> 
		sys_res_n	=> 
		
		calc_data	=> 
		calc_data2	=> 
		calc_operator	=> 
		calc_start	=> 
		calc_finished	=> 
		calc_result	=> 
		calc_status	=> 
		

	)
	
end architecture struct;
