-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.1 Build 222 10/21/2009 SJ Full Version
-- Created on Mon Apr 26 15:03:50 2010

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mjl_stratix_testSM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC
    );
END mjl_stratix_testSM;

ARCHITECTURE BEHAVIOR OF mjl_stratix_testSM IS
    TYPE type_fstate IS (state1,state2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
        ELSE
            CASE fstate IS
                WHEN state1 =>
                    reg_fstate <= state2;
                WHEN state2 =>
                    reg_fstate <= state1;
                WHEN OTHERS => 
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
